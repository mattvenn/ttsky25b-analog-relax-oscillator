magic
tech sky130A
magscale 1 2
timestamp 1762791078
<< psubdiff >>
rect 21282 6460 21306 7326
rect 22216 6460 22240 7326
<< psubdiffcont >>
rect 21306 6460 22216 7326
<< locali >>
rect 22500 9374 23340 9380
rect 21800 9317 22200 9320
rect 21800 9283 22163 9317
rect 22197 9283 22200 9317
rect 21800 9280 22200 9283
rect 22500 9226 23186 9374
rect 23334 9226 23340 9374
rect 22500 9220 23340 9226
rect 21290 6460 21306 7326
rect 22216 6460 22232 7326
<< viali >>
rect 12506 10806 12574 10874
rect 13826 10806 13894 10874
rect 22163 9283 22197 9317
rect 23186 9226 23334 9374
rect 5298 7818 5382 8040
rect 6610 7802 6698 8008
rect 19894 7906 19984 8132
rect 8926 7016 9088 7080
rect 17338 7018 17512 7088
<< metal1 >>
rect 4580 12520 21380 13400
rect 2820 12360 21380 12520
rect 2820 11620 2980 12360
rect 3901 12300 4059 12360
rect 4580 12000 21380 12360
rect 10760 11901 10840 12000
rect 3500 11780 4000 11800
rect 3500 11700 4080 11780
rect 3920 11680 4080 11700
rect 3920 11620 7080 11680
rect 3920 11520 6940 11620
rect 7040 11520 7080 11620
rect 8970 11650 9070 11656
rect 10760 11600 10841 11901
rect 4240 8000 4400 11520
rect 6940 11180 7040 11520
rect 8970 11150 9070 11550
rect 10300 11300 10841 11600
rect 11000 11400 11450 11500
rect 10760 11260 10841 11300
rect 8022 10900 8142 10906
rect 7180 10780 8022 10900
rect 8142 10780 8820 10900
rect 8022 10774 8142 10780
rect 5060 8040 6900 8080
rect 4240 7840 4860 8000
rect 2900 7300 3600 7500
rect 4240 7400 4400 7840
rect 5060 7818 5298 8040
rect 5382 8008 6900 8040
rect 5382 7818 6610 8008
rect 5060 7802 6610 7818
rect 6698 7802 6900 8008
rect 5060 7760 6900 7802
rect 3940 7240 4400 7400
rect 4240 6780 4400 7240
rect 4900 6780 5060 7240
rect 4240 6620 5060 6780
rect 5860 6140 6180 7760
rect 9150 7330 9900 7430
rect 8894 7080 9118 7098
rect 8894 7016 8926 7080
rect 9088 7016 9118 7080
rect 8894 6140 9118 7016
rect 9750 6450 9850 7330
rect 10400 6900 11100 7100
rect 11350 6850 11450 11400
rect 11660 11080 11740 12000
rect 11660 11000 12020 11080
rect 12500 10874 12580 12000
rect 12500 10806 12506 10874
rect 12574 10806 12580 10874
rect 12500 10794 12580 10806
rect 13820 10874 13900 12000
rect 14700 11080 14780 12000
rect 15560 11500 15640 12000
rect 16640 11994 16740 12000
rect 17344 11550 17350 11650
rect 17450 11550 17456 11650
rect 19550 11620 19650 11626
rect 15200 11200 15640 11500
rect 15800 11300 16350 11400
rect 15560 11160 15640 11200
rect 14380 11000 14780 11080
rect 13820 10806 13826 10874
rect 13894 10806 13900 10874
rect 13820 10794 13900 10806
rect 13564 9210 13570 9310
rect 13670 9210 13676 9310
rect 12790 8770 12890 8776
rect 12790 7490 12890 8670
rect 12350 7390 12890 7490
rect 12150 6860 12250 7210
rect 12790 6860 12890 7390
rect 13570 8214 13670 9210
rect 14320 8654 14560 8814
rect 13570 8054 13680 8214
rect 13570 7490 13670 8054
rect 13570 7390 14030 7490
rect 16250 7450 16350 11300
rect 17350 11170 17450 11550
rect 19550 11210 19650 11520
rect 18414 10920 18534 10926
rect 17560 10800 18414 10920
rect 18534 10800 19420 10920
rect 18414 10794 18534 10800
rect 20240 9880 20560 12000
rect 22480 11850 22580 11856
rect 23362 11850 24528 12186
rect 22580 11750 24528 11850
rect 22480 11744 22580 11750
rect 23362 11066 24528 11750
rect 20220 9560 22960 9880
rect 20920 9350 21060 9400
rect 23320 9380 24500 9800
rect 20920 9250 20930 9350
rect 21030 9320 21060 9350
rect 23174 9374 24500 9380
rect 22151 9320 22209 9323
rect 21030 9317 22209 9320
rect 21030 9283 22163 9317
rect 22197 9283 22209 9317
rect 21030 9280 22209 9283
rect 21030 9250 21060 9280
rect 22151 9277 22209 9280
rect 20920 9220 21060 9250
rect 23174 9226 23186 9374
rect 23334 9226 24500 9374
rect 23174 9220 24500 9226
rect 20200 8740 22940 9060
rect 20200 8180 20520 8740
rect 23320 8680 24500 9220
rect 19660 8132 20520 8180
rect 19660 7906 19894 8132
rect 19984 7906 20520 8132
rect 19660 7860 20520 7906
rect 16250 7430 16450 7450
rect 13570 6860 13670 7390
rect 16250 7350 17230 7430
rect 16300 7330 17230 7350
rect 14170 6860 14270 7160
rect 11500 6850 12900 6860
rect 11350 6760 12900 6850
rect 13560 6760 14900 6860
rect 15200 6800 15900 7100
rect 11350 6750 11750 6760
rect 11550 6450 11650 6750
rect 9750 6350 11650 6450
rect 14750 6450 14850 6760
rect 16350 6450 16450 7330
rect 14750 6350 16450 6450
rect 17286 7088 17586 7096
rect 17286 7018 17338 7088
rect 17512 7018 17586 7088
rect 17286 6140 17586 7018
rect 20200 6140 20520 7860
rect 21254 6140 22334 7462
rect 4280 5060 22334 6140
<< via1 >>
rect 6940 11520 7040 11620
rect 8970 11550 9070 11650
rect 8022 10780 8142 10900
rect 17350 11550 17450 11650
rect 13570 9210 13670 9310
rect 12790 8670 12890 8770
rect 19550 11520 19650 11620
rect 18414 10800 18534 10920
rect 22480 11750 22580 11850
rect 20930 9250 21030 9350
<< metal2 >>
rect 16470 11750 22480 11850
rect 22580 11750 22586 11850
rect 16470 11650 16570 11750
rect 17350 11650 17450 11656
rect 6940 11620 7040 11626
rect 7040 11520 7970 11620
rect 8070 11520 8079 11620
rect 8964 11550 8970 11650
rect 9070 11550 9970 11650
rect 6940 11514 7040 11520
rect 8016 10780 8022 10900
rect 8142 10780 8148 10900
rect 8022 4426 8142 10780
rect 9870 9310 9970 11550
rect 16470 11550 17350 11650
rect 18295 11620 18385 11624
rect 13570 9310 13670 9316
rect 9870 9210 13570 9310
rect 13570 9204 13670 9210
rect 16470 8770 16570 11550
rect 17350 11544 17450 11550
rect 18290 11615 19550 11620
rect 18290 11525 18295 11615
rect 18385 11525 19550 11615
rect 18290 11520 19550 11525
rect 19650 11520 19678 11620
rect 18295 11516 18385 11520
rect 20950 11418 21050 11750
rect 20930 11150 21050 11418
rect 18408 10800 18414 10920
rect 18534 10800 18540 10920
rect 12784 8670 12790 8770
rect 12890 8670 16570 8770
rect 18414 4742 18534 10800
rect 20930 9350 21030 11150
rect 20930 9244 21030 9250
rect 18414 4524 18536 4742
rect 18416 4447 18536 4524
rect 8022 4306 8732 4426
rect 8852 4306 8861 4426
rect 18412 4337 18421 4447
rect 18531 4337 18540 4447
rect 18416 4332 18536 4337
<< via2 >>
rect 7970 11520 8070 11620
rect 18295 11525 18385 11615
rect 8732 4306 8852 4426
rect 18421 4337 18531 4447
<< metal3 >>
rect 7965 11620 8075 11625
rect 7965 11520 7970 11620
rect 8070 11615 18390 11620
rect 8070 11525 18295 11615
rect 18385 11525 18390 11615
rect 8070 11520 18390 11525
rect 7965 11515 8075 11520
rect 18416 4447 18536 4452
rect 8727 4426 8857 4431
rect 8727 4306 8732 4426
rect 8852 4306 9046 4426
rect 9166 4306 9172 4426
rect 18416 4377 18421 4447
rect 18531 4377 18536 4447
rect 8727 4301 8857 4306
rect 18416 4259 18417 4377
rect 18535 4259 18536 4377
rect 18416 4258 18536 4259
rect 18417 4253 18535 4258
<< via3 >>
rect 9046 4306 9166 4426
rect 18417 4337 18421 4377
rect 18421 4337 18531 4377
rect 18531 4337 18535 4377
rect 18417 4259 18535 4337
<< metal4 >>
rect 17438 4484 19430 4588
rect 17438 4440 17542 4484
rect 9045 4426 9167 4427
rect 9668 4426 17542 4440
rect 9045 4306 9046 4426
rect 9166 4336 17542 4426
rect 19326 4440 19430 4484
rect 17718 4377 18536 4378
rect 9166 4306 9834 4336
rect 9045 4305 9167 4306
rect 9668 3884 9772 4306
rect 17718 4259 18417 4377
rect 18535 4259 18536 4377
rect 19326 4336 20330 4440
rect 17718 4258 18536 4259
rect 17718 4230 17838 4258
rect 16658 4226 17838 4230
rect 12932 4122 17838 4226
rect 12932 2934 13036 4122
rect 16658 4110 17838 4122
rect 16944 4000 17048 4110
rect 20226 2812 20330 4336
use sky130_fd_pr__res_high_po_0p69_QFH5ZW  sky130_fd_pr__res_high_po_0p69_QFH5ZW_0
timestamp 1762791078
transform 1 0 2935 0 1 9582
box -235 -2582 235 2582
use sky130_fd_pr__res_high_po_0p69_QFH5ZW  sky130_fd_pr__res_high_po_0p69_QFH5ZW_1
timestamp 1762791078
transform 1 0 10435 0 1 9182
box -235 -2582 235 2582
use sky130_fd_pr__res_high_po_0p69_QFH5ZW  sky130_fd_pr__res_high_po_0p69_QFH5ZW_2
timestamp 1762791078
transform 1 0 3535 0 1 9582
box -235 -2582 235 2582
use sky130_fd_pr__res_high_po_0p69_QFH5ZW  sky130_fd_pr__res_high_po_0p69_QFH5ZW_3
timestamp 1762791078
transform 1 0 15835 0 1 9182
box -235 -2582 235 2582
use sky130_fd_pr__res_high_po_0p69_QFH5ZW  sky130_fd_pr__res_high_po_0p69_QFH5ZW_4
timestamp 1762791078
transform 1 0 11035 0 1 9182
box -235 -2582 235 2582
use sky130_fd_pr__res_high_po_0p69_QFH5ZW  sky130_fd_pr__res_high_po_0p69_QFH5ZW_5
timestamp 1762791078
transform 1 0 15235 0 1 9182
box -235 -2582 235 2582
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1704896540
transform 1 0 21386 0 1 9068
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_8  x1
timestamp 1704896540
transform 1 0 21478 0 1 9068
box -38 -48 1234 592
use sky130_fd_pr__cap_mim_m3_1_39BNLG  XC1
timestamp 1710760421
transform 1 0 9866 0 1 -11812
box -3186 -15800 3186 15800
use sky130_fd_pr__cap_mim_m3_1_39BNLG  XC2
timestamp 1710760421
transform 1 0 17142 0 1 -11696
box -3186 -15800 3186 15800
use sky130_fd_pr__nfet_01v8_L9BG78  XM1
timestamp 1710760421
transform 1 0 8996 0 1 9210
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_L9BG78  XM2
timestamp 1710760421
transform 1 0 17396 0 1 9210
box -396 -2210 396 2210
use sky130_fd_pr__pfet_01v8_5Q5MA6  XM3
timestamp 1710760421
transform 1 0 14196 0 1 9219
box -396 -2219 396 2219
use sky130_fd_pr__pfet_01v8_5Q5MA6  XM4
timestamp 1710760421
transform 1 0 12196 0 1 9219
box -396 -2219 396 2219
use sky130_fd_pr__nfet_01v8_L9BG78  XM5
timestamp 1710760421
transform 1 0 4996 0 1 9210
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_L9BG78  XM6
timestamp 1710760421
transform 1 0 6996 0 1 9210
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_L9BG78  XM8
timestamp 1710760421
transform 1 0 19596 0 1 9210
box -396 -2210 396 2210
<< labels >>
flabel metal1 5140 12500 5340 12700 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 4660 5360 4860 5560 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 23380 9240 23580 9440 0 FreeSans 256 0 0 0 osc_out
port 2 nsew
flabel metal1 12790 6760 12890 8670 0 FreeSans 1600 0 0 0 osc_a
flabel metal1 13570 6760 13670 9210 0 FreeSans 1600 0 0 0 osc_b
flabel metal2 8022 4306 8142 10780 0 FreeSans 1600 0 0 0 left_cap
flabel space 18414 4230 18534 10800 0 FreeSans 1600 0 0 0 right_cap
flabel metal1 4240 11520 6940 11680 0 FreeSans 1600 0 0 0 cset
flabel metal1 23362 11066 24528 12186 0 FreeSans 1600 0 0 0 osc_a
port 3 nsew
<< end >>
